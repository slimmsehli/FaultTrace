
package i2c_package;

`include "uvm_macros.svh"
import uvm_pkg::*;

`include "i2c_item.sv"
`include "i2c_driver.sv"
`include "i2c_agent.sv"
`include "i2c_sequences.sv"
`include "i2c_tests.sv"

endpackage
